library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY RAM_1P_16N_8N is
		generic(BitsOfAddress  : natural := 4;
				  BitsInDataOfAddress : natural := 8);
				  
		port(Clk : in std_logic;
			  Enable : in std_logic;
			  writeData : in std_logic_vector(BitsInDataOfAddress -1 downto 0);--wite on 8bits of case x"XX"
			  address : in std_logic_vector(BitsOfAddress-1 downto 0); --cases 16
			  readData : out std_logic_vector(BitsInDataOfAddress -1 downto 0)); --read the 8 bits

end RAM_1P_16N_8N;

architecture Behavioral of RAM_1P_16N_8N is
subtype TDataWord is std_logic_vector(BitsInDataOfAddress -1 downto 0);
type TMemory is array (0 to 2*BitsOfAddress -1) of TDataWord;
signal s_memory : TMemory;
begin
	process(Clk)
			begin
					if(rising_edge(Clk))then
						if (Enable = '1') then
							s_memory(to_integer(unsigned(address))) <= writeData;
						end if;
					end if;
			end process;
			readData <= s_memory(to_integer(unsigned(address)));
end Behavioral;			  